module vz32_decoder()

endmodule

module regfile_32x32()

endmodule

module regfile_16x64()

endmodule

module alu()

endmodule

module fp()

endmodule

module vz32_plain()

endmodule